// barrel shifter 

module barrel_shifter(operand2, cin); 
    
endmodule
